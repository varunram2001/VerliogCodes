module xnor_gate(c,a,b);
input a,b;
output c;
xnor (c,a,b);
endmodule
