module testbench;

  reg clk;
  reg reset;
  wire [3:0] count;

  johnson_counter uut (
    .clk(clk),
    .reset(reset),
    .count(count)
  );

  initial begin
    // Open VCD file for waveform dumping
    $dumpfile("waveform.vcd");
    $dumpvars(0, testbench); // Dump all variables
    
    // Initialize inputs
    clk = 0;
    reset = 0;
    
    // Apply inputs and check outputs
    #5 reset = 1;
    #5 reset = 0;
    #10 clk = 1; #5 clk = 0; // Shift counter (0001 -> 1000)
    #10 clk = 1; #5 clk = 0; // Shift counter (1000 -> 1100)
    #10 clk = 1; #5 clk = 0; // Shift counter (1100 -> 1110)
    #10 clk = 1; #5 clk = 0; // Shift counter (1110 -> 1111)
    #10 clk = 1; #5 clk = 0; // Shift counter (1111 -> 0111)
    #10 clk = 1; #5 clk = 0; // Shift counter (0111 -> 0011)
    #10 clk = 1; #5 clk = 0; // Shift counter (0011 -> 0001)
    #10 clk = 1; #5 clk = 0; // Shift counter (0001 -> 1000)
    
    // Finish simulation
    $finish;
  end

endmodule
