// Code your design here
//OR gate using Structural modeling
module or_gate_s(a,b,y);
input a,b;
output y;

or(y,a,b);
                
endmodule